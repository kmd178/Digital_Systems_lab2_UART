`timescale 1ns / 1ps
module systemUART(
    );


endmodule
